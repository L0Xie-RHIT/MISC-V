module Control(
    input [2:0] opcode,
    input [3:0] func,
    input reset,
    output reg RegWrite,
    output reg ALUSrc,
    output reg [2:0] ALUOp,
    output reg RegStore,
    output reg MemWrite,
    output reg MemRead,
    output reg Branch
);


endmodule